/****************************************************************************
 * uvm_sdv_memblk_connector_pkg.sv
 ****************************************************************************/

/**
 * Package: uvm_sdv_memblk_connector_pkg
 * 
 * TODO: Add package documentation
 */
`include "uvm_macros.svh"
package uvm_sdv_memblk_connector_pkg;
	import uvm_sdv_pkg::*;
	
	`include "memblk_connector/uvm_sdv_memblk_connector.svh"
endpackage


