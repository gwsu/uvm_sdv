
`include "uvm_macros.svh"
package types_pkg;
	import uvm_pkg::*;
	
	`include "sw_txn.svh"
	`include "sw_txn_seq.svh"
	`include "sw_txn_driver.svh"
	
endpackage

