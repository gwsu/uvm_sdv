
`include "uvm_macros.svh"

package simple_dpi_env_pkg;
	import uvm_pkg::*;
	import uvm_sdv_pkg::*;
	import uvm_sdv_dpi_pkg::*;
	import types_pkg::*;

	`include "simple_dpi_sdv_connector.svh"
	`include "simple_dpi_env.svh"
	
endpackage
