/****************************************************************************
 * uvm_sdv_agent_if.svh
 ****************************************************************************/
`ifndef INCLUDED_uvm_sdv_agent_if_svh
`define INCLUDED_uvm_sdv_agent_if_svh

/**
 * Class: uvm_sdv_agent_if
 * 
 * TODO: Add class documentation
 */
virtual class uvm_sdv_agent_if;
	
	virtual task queue_msg();
	endtask

endclass

`endif /* INCLUDED_uvm_sdv_agent_if_svh */
